module RGB_Overwrite(
input [10:0] vga_x,vga_y,
input clk,
output [7:0] box_r,
output [7:0] box_g,
output [7:0] box_b
);


//always @(*) begin
//	if (inBox1) begin
//		box_r = 244;
//		box_g = 214;
//		box_b = 158;
//	end
////	else if(inBox1) begin
////		box_r = 10;
////		box_g = 10;
////		box_b = 10;
////	end
//	else
//		box_r = 0;
//		box_g = 0;
//		box_b = 0;
//end

endmodule 