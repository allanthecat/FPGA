module Line_Buffer_3_Taps(
input clk,
input en,
input [7:0] grey_in,
output [7:0] r0,r1,r2
);




endmodule 